`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   16:22:39 09/06/2021
// Design Name:   MEMORY_V
// Module Name:   C:/Users/donal/Documents/adld/bram_attempt_4/drtb.v
// Project Name:  bram_attempt_4
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: MEMORY_V
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module drtb;

	// Inputs
	reg clka;
	reg [5:0] address;

	// Outputs
	wire [19:0] douta;

	// Instantiate the Unit Under Test (UUT)
	MEMORY_V uut (
		.clka(clka), 
		.address(address), 
		.douta(douta)
	);

	initial begin
		// Initialize Inputs
		clka = 0;
		address = 0;

		// Wait 100 ns for global reset to finish
		#1;
        
		// Add stimulus here
		clka = 0;
		address = 0;
		#3;
		clka=1;
		#1;
		#1;
        
		// Add stimulus here
		clka = 0;
		address = 1;
		#3;
		clka=1;
		#1;
		#1;
        
		// Add stimulus here
		clka = 0;
		address = 2;
		#3;
		clka=1;
		#1;
		
		clka = 0;
		address = 3;
		#3;
		clka=1;
		#1;
		
		clka = 0;
		address = 4;
		#3;
		clka=1;
		#1;
		
		
		clka = 0;
		address = 5;
		#3;
		clka=1;
		#1;
		
		
		clka = 0;
		address = 6;
		#3;
		clka=1;
		#1;
		
		
		clka = 0;
		address = 2;
		#3;
		clka=1;
		#1;
		
		
		clka = 0;
		address = 2;
		#3;
		clka=1;
		#1;
		
		
		clka = 0;
		address = 2;
		#3;
		clka=1;
		#1;

	end
      
endmodule

