`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:15:45 09/06/2021 
// Design Name: 
// Module Name:    MEMORY_V 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module working_clk(
	input clk,
	output reg clock,
	output reg clk1
	);
	reg [24:0] counter;
	initial counter=5'b0;
	always @(posedge clk) begin
		counter<=counter +1'b1;
		if (counter[4:0]==5'b0)
			clock<=1'b1;
		else begin
			if (counter[4:0]==5'b1)
				clock<=1'b0;
			end
		if (counter==25'b0)
			clk1<=1'b1;
		else begin
			if (counter==25'b1)
				clk1<=1'b0;
			end
		end
	endmodule

module MEMORY_V(
    input clka,
    output wire [19:0] douta,
	 output wire clock,
	 output wire clk1,
	 output reg [1:0] X,
	 output reg [6:0] Y,
	 output reg [1:0] D,
	 output reg [5:0] address
    );
	reg [7:0] mem [15:0];
	initial address=6'b0;
	reg [7:0] A;
	reg [7:0] B;
	reg [7:0] x;
	reg [3:0] R;
	reg count2 =1'b0;
	
	working_clk random(clka,clock,clk1);
	mem temp(.clka(clock),.addra(address),.douta(douta));
	
	always @(posedge clk1) begin
		case (douta[19:16])
		1:	begin
			A=mem[douta[15:12]];
			B=mem[douta[11:8]];
			case(douta[3:0])
				0: mem[douta[7:4]]=A;
				1: {D[1],mem[douta[7:4]]}= (~A+9'b1);
				2: {D[1],mem[douta[7:4]]}= A+B+9'b0;
				3: {D[1],mem[douta[7:4]]}=A+(9'b1+(~B));
				4: {D[1],mem[douta[7:4]]}= (A+9'b00000)<<1;
				5: {D[1],mem[douta[7:4]]}= (A+9'b00000)>>1;
				6: {D[1],mem[douta[7:4]]}=A+9'b1;
				7: begin
					mem[douta[7:4]]=A-8'b1;
					if (A<1)
						D[1]=1;
					end
				8: mem[douta[7:4]]=~A;
				9: mem[douta[7:4]]=A&B;
				10: mem[douta[7:4]]=A|B;
				11: mem[douta[7:4]]=A^B;
				12: mem[douta[7:4]]=A<<1;
				13: mem[douta[7:4]]=A>>1;
				14: mem[douta[7:4]]=A;
				15: mem[douta[7:4]]=8'b11111111;
				endcase
				if(mem[douta[7:4]]==8'b0)
					D[0]=1;
				x=mem[douta[7:4]];
			end
		4: begin
			address=address+douta[5:0];
			end
		7: begin
			if (D[0]) begin
				address=address+douta[5:0];
				end
			end
		5:	begin
			if (D[1])
				address=address+douta[5:0];
			end
		6:	begin
			if (D[1]==0)
				address=address+douta[5:0];
			end
		endcase
		address=address+1'b1;
		end
				
	always @(posedge clock) begin
		X={X[0],X[1]};
		case(count2)
			0:R=x[3:0];
			1:R=x[7:4];
		endcase
		count2=count2+1'b1;
		end
	
	always @(R)
			begin
			case(R)
			0:Y=7'b0000001;
			1:Y=7'b1001111;
			2:Y=7'b0010010;
			3:Y=7'b0000110;
			4:Y=7'b1001100;
			5:Y=7'b0100100;
			6:Y=7'b0100000;
			7:Y=7'b0001111;
			8:Y=7'b0000000;
			9:Y=7'b0001100;
			10:Y=7'b0001000;
			11:Y=7'b1100000;
			12:Y=7'b0110001;
			13:Y=7'b1000010;
			14:Y=7'b0110000;
			15:Y=7'b0111000;
			default: Y=7'b1111111;
			endcase
			end
endmodule
