//`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    02:04:56 07/29/2021 
// Design Name: 
// Module Name:    dancing_lights 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module dancing_lights(
    input clk,
    input reset,
    output reg [23:0]ctr,
    output reg working_clk=0,
    output reg [3:0] x,
    output reg [7:0] y
    );
always@ (posedge  clk)
begin
  if (reset)
  begin 
	 ctr <= 24'b0;
  end
  else
  begin
     if (ctr == 24'b1)
	  begin 
	   ctr <= 24'b0;
	end
	else
	begin
	ctr <= ctr + 1'b1;
	end
  end
 end
 always @(posedge ctr[23])
 begin 
 if (reset) begin
 y = 8'b11111110;
 x = 4'b110;
 end
 else
 begin
 if (y == 8'b01111111) begin
 x = ((x<<1) | (x>>3));
 end
 y = ((y<<1) | (y>>7));

end 
end

endmodule
	 
